library ieee;
use ieee.std_logic_1164.all;

entity one_pulse is
	port (
		clk		: in std_ulogic;
		rst		: in std_ulogic;
		input	: in std_ulogic;
		pulse	: out std_ulogic);
end entity;

architecture one_pulse_arch of one_pulse is
	
	begin
	
end architecture;
